library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fixed_mult is
    generic ( WIDTH : integer := 16 );
    port (
        a, b : in std_logic_vector(WIDTH-1 downto 0);
        result : out std_logic_vector(WIDTH-1 downto 0)
    );
end fixed_mult;

architecture rtl of fixed_mult is
begin
    process(a, b)
        variable v_a, v_b : signed(WIDTH-1 downto 0);
        variable v_res_full : signed(2*WIDTH-1 downto 0);
    begin
        v_a := signed(a);
        v_b := signed(b);
        v_res_full := v_a * v_b;
        
        -- Q1.15 * Q1.15 = Q2.30
        -- ????? ????? ????? ?? ????? Q1.15.
        -- ??? ?????? ?? ?????? ???????? (??????? ?? ?-LSB ???????? ??? ??? ????? ?????)
        -- ???? ??? ?????? ?? 30 downto 15
        result <= std_logic_vector(v_res_full(WIDTH + WIDTH - 2 downto WIDTH - 1));
    end process;
end rtl;
